module vrobot

/*
struct C.INPUT

pub fn type_stuff() {
  // Keyboard
  input := &C.INPUT{}
  vkey := C.VK_RETURN
  input.type = 1 // C.INPUT_KEYBOARD
  input.ki.wScan = C.MapVirtualKey(vkey, C.MAPVK_VK_TO_VSC)
  input.ki.time = 0 
  input.ki.dwExtraInfo = 0
  input.ki.wVk = vkey
  input.ki.dwFlags = 0
  C.SendInput(1, &input, sizeof(C.INPUT))

  input.ki.dwFlags = C.KEYEVENTF_KEYUP
  C.SendInput(1, &input, sizeof(C.INPUT))
}
*/
